library IEEE;
use IEEE.std_logic_1164.all;

entity neander_rom is
	port (
		mclk: in std_logic;
		btn: in std_logic_vector(3 downto 0);
		a_to_g: out std_logic_vector (6 downto 0);
		an: out std_logic_vector(3 downto 0);
		dp: out std_logic
	);
end neander_rom;

architecture neander_rom of neander_rom is
component x7seg
	port (
		x: in std_logic_vector(15 downto 0);
		clk: in std_logic ;
		clr: in std_logic ;
		a_to_g: out	std_logic_vector (6 downto 0);
		an:     out std_logic_vector (3 downto 0);
		dp: out std_logic 
	);
end component;
component rom
	port (
		addr: in std_logic_vector (3 downto 0);
		M: out std_logic_vector (7 downto 0)
	);
end component;

signal memory_address: std_logic_vector (3 downto 0);
signal memory_output: std_logic_vector (7 downto 0);
begin
   memory_address <= not btn;

	U1: rom port map(
		addr => memory_address,
		M => memory_output
	);
	U2: x7seg port map (
		x => X"00" & memory_output,
		clk => mclk,
		clr => '0',
		a_to_g => a_to_g,
		an => an,
		dp => dp
	);


end neander_rom;